package timer_pkg;

`include "packet.sv"
`include "stimulus.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "environment.sv"

endpackage